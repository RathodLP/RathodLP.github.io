module top;

initial begin
	$display("Welcome to GitHub");
	$display("Write SV Code");
	$display("Hi Rathod");
end
endmodule
