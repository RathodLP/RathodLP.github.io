> Hi This is sample file for SV
> #Hello world
